module case_theoretical;

    // case, casex, casez
    // case - all the bits must be exactly same
    // casex - not considering x, z values
    // casez - not considering z's

    case (expression)
        case_item0: statement_1;
        case_item2: statement_2;
        default: statement_default;
    endcase

endmodule