module short_long_int_integer_example;

    // 16 - bit signed integer - 2 bytes
    // -32768 until 32767
    /* 
    32,767 → Binary: 01111111 11111111.
    -32,768 → Binary: 10000000 00000000.

    Operations:
    Arithmetic: +, -, *, /, %.
    Bitwise: &, |, ^, ~.
    Shift: <<, >>, >>>.
    Comparison: <, <=, >, >=, ==, !=.
    */


    // 64 - bits - signed integer - 8 bytes
    // Range: -9,223,372,036,854,775,808 to 9,223,372,036,854,775,807 (signed).

    /* 
    9,223,372,036,854,775,807 → Binary:
    01111111 11111111 11111111 11111111 11111111 11111111 11111111 11111111

    -9,223,372,036,854,775,807 → Binary:
    10000000 00000000 00000000 00000000 00000000 00000000 00000000 00000001
    */

    // Integer - Int


endmodule