module dynamic_array;




endmodule
