module while_concept;




endmodule